module test_bench;
endmodule