module test ();
endmodule