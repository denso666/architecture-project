`timescale 1ns/1ns
module and1b ( input A, B, output R );

    assign R = A & B;

endmodule // and
