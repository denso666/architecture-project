module buffer_wb (
    input clk,
    input [1:0] in,
    output reg [1:0] out
);

    always @ (posedge clk) begin
        out = in;
    end

endmodule // buffer_wb
